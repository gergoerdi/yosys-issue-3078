module Top(
           output [5:2] LED
           );

   assign LED[5:2] = 4'b1101;
   
endmodule
